library	ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;   

entity ROM is
	port(	addr		: in std_logic_vector(15 downto 0);
			data_out	: out std_logic_vector(15 downto 0));
end entity;

architecture struct of ROM is

type mem_type is array (0 to 31) of std_logic_vector(15 downto 0);
/*signal mem: mem_type:=(	0 => "0001100100111111",	--ADI R4 R4 11111   		
								1 => "0001101101001111",	--ADI R5 R5 00010	
								2 => "0111110000110000",	--SM R6 00110000
								3 => "0101100110000001",	--SW R4 R6 01	
								4 => "0011100000000000",	--LHI R4 0000
								5 => "0011101000000000",	--LHI R5 0000
								6 => "0001011011000111",	--ADI R3 R3 7

								7 => "0110101000000110",	--LM R5 00000110		
								
								8 => "1100001101000011",	--BEQ R1 R5 3
								9 => "0001001001111111",	--ADI R1 R1 -1
								10 => "1000110111111110",	--JAL R6 -2
								
								11 => "1100010101000100",	--BEQ R2 R5 4
								12=> "0001010010111111",	--ADI R2 R2 -1
								13=> "0100001101000001",	--LW R1 R5 1
								14=> "1000110111111010",	--JAL R6 -6
								
								15=> "0001000000000001",	--ADI R0 R0 1
								16=> "0000101011111000",	--JLR R6 R3
					
								others => "0000000000000000");*/

signal mem: mem_type:=(	0 => "0001100100000111",	--ADI R4 R4 11111   		
								1 => "0001101101000010",	--ADI R5 R5 00010	
								2 => "0111110000100000",	--SM R6 00100000
								3 => "0101100110000001",	--SW R4 R6 01	
								4 => "0011100000000000",	--LHI R4 0000
								5 => "0011101000000000",	--LHI R5 0000
								6 => "0001011011000111",	--ADI R3 R3 7

								7 => "0110101000000110",	--LM R5 00000110		
								
								8 => "1100001101000011",	--BEQ R1 R5 3
								9 => "0001001001111111",	--ADI R1 R1 -1
								10 => "1000110111111110",	--JAL R6 -2
								
								11 => "1100010101000100",	--BEQ R2 R5 4
								12=> "0001010010111111",	--ADI R2 R2 -1
								13=> "0100001101000001",	--LW R1 R5 1
								14=> "1000110111111010",	--JAL R6 -6
								
								15=> "0001000000000001",	--ADI R0 R0 1
								16=> "0011110000000000",	--LHI R6 0
								17=> "0001110110000011",	--ADI R6 R6 111111
								18=> "1100000110000010",	--BEQ R6 R0 +2
								19=> "0000101011111000",	--ADD R5 R3 R7
								20=> "0011000000000000",	--LHI R0 0
								21=> "0000101011111000",	--ADD R5 R3 R7
								others => "0000000000000000");	
		
/*signal mem: mem_type:=(	0 => "0001010010000010",	--ADI R2 R2 00010   		
								1 => "0001001001000010",	--ADI R1 R1 00010	
								
								2 => "1100001101000011",	--BEQ R1 R5 3
								3 => "0001001001111111",	--ADI R1 R1 -1
								4 => "1000110111111110",	--JAL R6 -2
								
								5 => "1100010101000100",	--BEQ R2 R5 4
								6 => "0001010010111111",	--ADI R2 R2 -1
								7 => "0001001001000010",	--ADI R1 R1 00010	
								8 => "1000110111111010",	--JAL R6 -6
								
								9 => "0001000000000001",	--ADI R0 R0 1
								10=> "1000110111110110",	--JAL R6 -10
					
								others => "0000000000000000");*/		
								
begin
	
	data_out <= mem(conv_integer(addr(4 downto 0)));
	
end struct;
